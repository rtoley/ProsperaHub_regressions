tests_cmp.sv