tests_modular.sv