tests_red.sv